module cache_control (
);

endmodule : cache_control

module cache #(
    parameter s_offset = 5,
    parameter s_index  = 3,
    parameter s_tag    = 32 - s_offset - s_index,
    parameter s_mask   = 2**s_offset,
    parameter s_line   = 8*s_mask,
    parameter num_sets = 2**s_index
)
(
);

cache_control control
(
);

cache_datapath datapath
(
);

bus_adapter bus_adapter
(
);

endmodule : cache
